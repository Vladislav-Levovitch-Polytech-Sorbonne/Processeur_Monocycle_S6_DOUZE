library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use IEEE.std_logic_unsigned.ALL;

entity test_bench_UAL_Banc_de_Registre_entity is
    
end test_bench_UAL_Banc_de_Registre_entity;

architecture test_bench_UAL_Banc_de_Registre_architecture of test_bench_UAL_Banc_de_Registre_entity is
	
	-- Entrees
	signal SIGNAL_Test_Bench_Clk_BRUAL, SIGNAL_Test_Bench_Rst_BRUAL, SIGNAL_Test_Bench_WE_BRUAL : std_logic := '0';
	signal SIGNAL_Test_Bench_Ra_BRUAL, SIGNAL_Test_Bench_Rb_BRUAL, SIGNAL_Test_Bench_Rw_BRUAL : std_logic_vector(3 downto 0) := "0000"; -- Bus Adresse
	signal SIGNAL_Test_Bench_OP_BRUAL  : std_logic_vector (2 downto 0) := "000"; -- 3 bits de Commande de l operation a selectionner sur l UAL
	
	-- Sorties
	signal SIGNAL_Test_Bench_N_BRUAL, SIGNAL_Test_Bench_Z_BRUAL, SIGNAL_Test_Bench_C_BRUAL, SIGNAL_Test_Bench_V_BRUAL : std_logic := '0'; -- Drapeaux
	signal SIGNAL_Test_Bench_S_BRUAL : std_logic_vector(31 downto 0) := x"0000_0000"; -- Bit de resultat

begin 


	UUT_UAL_Banc_de_Registre : entity work.UAL_Banc_de_Registre_entity
        port map 
		(

			Clk_BRUAL => SIGNAL_Test_Bench_Clk_BRUAL, 
			Rst_BRUAL => SIGNAL_Test_Bench_Rst_BRUAL, 
			WE_BRUAL  => SIGNAL_Test_Bench_WE_BRUAL,

			Ra_BRUAL => SIGNAL_Test_Bench_Ra_BRUAL,
			Rb_BRUAL => SIGNAL_Test_Bench_Rb_BRUAL,
			Rw_BRUAL => SIGNAL_Test_Bench_Rw_BRUAL,
			OP_BRUAL => SIGNAL_Test_Bench_OP_BRUAL,

			S_BRUAL => SIGNAL_Test_Bench_S_BRUAL,
			N_BRUAL => SIGNAL_Test_Bench_N_BRUAL, 
			Z_BRUAL => SIGNAL_Test_Bench_Z_BRUAL, 
			C_BRUAL => SIGNAL_Test_Bench_C_BRUAL,
			V_BRUAL => SIGNAL_Test_Bench_V_BRUAL
        );

	UUT_THE_HORLOGE : entity work.Tic_Tac_entity -- Horloge principale
        port map 
		(
            THE_Clk => SIGNAL_Test_Bench_Clk_BRUAL
        );

Test_bench_UAL_Banc_de_Registre : process 
	
    begin		

		-- Valeur initiale d entree
		wait for 1 ns; 
		SIGNAL_Test_Bench_WE_BRUAL <= '1';
		SIGNAL_Test_Bench_Rst_BRUAL <= '0'; -- Par securite 

		SIGNAL_Test_Bench_S_BRUAL <= x"0020_4010"; -- Valeur initiale pour R15
		SIGNAL_Test_Bench_Rw_BRUAL <= "1111"; -- R15
		wait for 12 ns;

		-- R(1) = R(15)
		SIGNAL_Test_Bench_Ra_BRUAL <= "1111"; -- R15
		wait for 1 ns; -- Meilleur lisibilite chronogramme
		SIGNAL_Test_Bench_OP_BRUAL <= "011";
		wait for 12 ns;

		wait;
    end process Test_bench_UAL_Banc_de_Registre;   
end test_bench_UAL_Banc_de_Registre_architecture;