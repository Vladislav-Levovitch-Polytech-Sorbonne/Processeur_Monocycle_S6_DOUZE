library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use IEEE.std_logic_unsigned.ALL; -- Pas super utile vu que numeric a deja et les signed et le unsigned mais par precaution pour eviter les bug on laisse

entity UAL_Unite_Arithmetique_et_Logique_TEST_BENCH_entity is
    port 
    (
        -- Test Bench
    );
end entity UAL_Unite_Arithmetique_et_Logique_TEST_BENCH_entity;

architecture UAL_Unite_Arithmetique_et_Logique_TEST_BENCH_architecture of UAL_Unite_Arithmetique_et_Logique_TEST_BENCH_entity is 

end architecture